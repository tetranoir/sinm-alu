module testbench();
// Declare inputs as regs and outputs as wires
reg [7:0] newpc;
reg clk;
reg wenable;
reg reset;


wire [7:0] currentpc;

// Initialize all variables
initial begin        
	clk = 1;       // initial value of clock
	reset = 0;  	// initial value of reset
	wenable = 0;     // initial value of wenable
	
	newpc = 2;      // initial value of newpc



	#10  reset = 1;    // use reset to set pc to 0
	#10  reset = 0;    // end of reset pulse.
	#10      // wait a cycle, make sure the PC doesn't change
	#10  wenable = 1; newpc = 4;    // set wenable high, pc should change
	#10  newpc = 5;   // try a few PC values
	#10  newpc = 7; 
	#10  reset = 1;   //see if reset works when wenable high
	#10  reset = 0; wenable = 0;

 end


// Clock generator
always begin
   #5  clk = ~clk; // Toggle clock every 5 ticks
						// this makes the clock cycle 10 ticks
end

// the following creates an instance of our program_counter register.
//   I copied this code verbatim from the walkthough.v that was
//   generated by Quartus when I created the .v file from the .bdf.

program_counter	b2v_inst(
	.clock(clk),
	.wenable_i(wenable),
	.reset_i(reset),
	.newpc_i(newpc),
	.pc_o(currentpc));


endmodule
